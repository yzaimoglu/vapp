module api