module controllers